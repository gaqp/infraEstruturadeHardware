module Mips(input clock);

endmodule 