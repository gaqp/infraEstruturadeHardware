module Mux_2_1();
endmodule 